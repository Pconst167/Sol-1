package pa_fpu;

  typedef enum logic[3:0]{
    op_add = 4'h0,
    op_sub = 4'h1,
    op_mul,
    op_square,
    op_div,
    op_sqrt,
    op_sin,
    op_cos,
    op_tan,
    op_ln,
    op_exp
  } e_fpu_operation;

  typedef enum logic[3:0]{
    arith_idle_st,
    arith_add_st,
    arith_sub_st,
    arith_mul_wait_st,
    arith_div_wait_st,

    arith_result_valid_st
  } e_arith_state;

  typedef enum logic [2:0]{
    mul_start_st,
    mul_product_add_st,
    mul_product_shift_st,
    mul_result_set_st,
    mul_end_st
  } e_mul_state;

  typedef enum logic[3:0]{
    main_idle_st,
    main_wait_st,
    main_finish_st,
    main_wait_ack_st,

    main_mul_wait_st
  } e_main_state;


endpackage